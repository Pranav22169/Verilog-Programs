module decoder3to8(E, i0, i1, i2, y0, y1, y2, y3, y4, y5, y6, y7);
input E, i0, i1, i2; 
output y0, y1, y2, y3, y4, y5, y6, y7;
reg y0, y1, y2, y3, y4, y5, y6, y7; 

always @*
begin 
    

